`include "../01_RTL/IOTDF.v"
`include "../01_RTL/crc_sort_core.v"
`include "../01_RTL/des_core.v"