// list all paths to your design files
`include "../01_RTL/core.v"
`include "../01_RTL/conv_3x3.v"
`include "../sram_512x8/sram_512x8.v"

